#! COINCIDENCE Circuit.

* A COINCIDENCE gate is supposed to fire only if its inputs arrive simultaneously.
* For its implementation, we use an RSFQ AND gate.


* Testbench
.tran 1p 0.8n
.options ysep
R10 10 11 100
R11 20 21 100
R12 30 31 100
V0 VCC 0 pwl 0 0 10p 10m

* Input Logic Pulses
V1 10 0 pulse 0 50m 200p 50p 50p 100p 350p
V2 20 0 pulse 0 50m 100p 50p 50p 100p 700p

* Reset Pulse / Clock
V3 30 0 pulse 0 50m 10p 50p 50p 100p 300p

* Macroscopic Coincidence Circuit
X0 11 12 VCC dcsfq
X1 12 IN1 VCC jtl

X2 21 22 VCC dcsfq
X3 22 IN2 VCC jtl

X4 31 CLK VCC dcsfq

X7 IN1 IN2 CLK OUT VCC cin


* RSFQ Pulse Generation
* RS = JJ damping shunts, using Stewart-McCumber parameter with B_c = 1
.subckt dcsfq IN OUT VBIAS
B0 9 5 15 jjr ics=170uA
RS0 9 5 4
B1 10 11 16 jjr ics=250uA
RS1 10 11 2.7
B2 12 13 17 jjr ics=150uA
RS2 12 13 4.6
B3 7 14 18 jjr ics=170uA
RS3 7 14 4

L0 12 0 3.58pH
LP0 8 6 0.08pH
LP1 4 9 1.29pH
LP2 5 6 1.13pH
LP3 6 10 1.74pH
LP4 5 7 0.21pH
LP5 4 12 1.27pH
LP6 11 0 0.13pH
LP7 13 7 0.69pH
LP8 14 0 0.18pH

LT0 10 OUT 2.11pH
LT1 IN 4 3.38pH

R0 VBIAS 8 27
.ends dcsfq



* Single JTL Circuit Element
.subckt jtl IN OUT VBIAS
B0 5 7 9 jjr ics=250uA
RS0 5 7 2.7
B1 6 8 10 jjr ics=250uA
RS1 6 8 2.7

LP0 7 0 .1pH
LP1 8 0 .1pH

LT0 IN 5 2.1pH
LT1 5 4 2.1pH
LT2 4 6 2.1pH
LT3 6 OUT 2.1pH

R0 VBIAS 4 29
.ends jtl

* Single JTL Circuit Element for pseudo-"level shifting" to lower Ic
.subckt jtl_lo IN OUT VBIAS
B0 5 7 9 jjr ics=150uA
RS0 5 7 4.6
B1 6 8 10 jjr ics=150uA
RS1 6 8 4.6

LP0 7 0 .1pH
LP1 8 0 .1pH

LT0 IN 5 3.5pH
LT1 5 4 3.5pH
LT2 4 6 3.5pH
LT3 6 OUT 3.5pH

R0 VBIAS 4 30
.ends jtl_lo


* Splitter Element
.subckt split IN OUT1 OUT2 VBIAS
B0 2 0 100 jjr ics=355uA
R0 2 0 1.9
B1 7 0 101 jjr ics=250uA
R2 7 0 2.7
B2 9 0 102 jjr ics=250uA
R3 9 0 2.7

L0 IN 1 0.8p
L1 1 3 1.2p
L2 3 5 0.05p
L3 5 6 1.6p
L4 6 OUT1 1.98p
L5 5 8 1.6p
L6 8 OUT2 1.98p

LP0 1 2 0.05p
LP1 4 3 0.13p
LP2 6 7 0.05p
LP3 8 9 0.05p

R1 VBIAS 4 16.7
.ends split


* Single Coincidence Element
.subckt cin IN1 IN2 CLK OUT VBIAS
* Clock signal is 
X5 CLK CLK1 CLK2 VBIAS split

L0 IN1 40 2p
L1 41 43 10p
L2 CLK1 42 2p
L3 43 47 4p
L4 IN2 50 2p
L5 44 46 10p
L6 CLK2 45 2p
L7 46 48 4p
L8 49 OUT 1.5p

B0 40 41 100 jjr ics=175uA
B1 41 0 101 jjr ics=175uA
B2 43 0 102 jjr ics=250uA
B3 42 43 103 jjr ics=175uA
B4 47 49 104 jjr ics=175uA
B5 50 44 105 jjr ics=175uA
B6 44 0 106 jjr ics=175uA
B7 46 0 107 jjr ics=250uA
B8 45 46 108 jjr ics=175uA
B9 48 49 109 jjr ics=175uA
B10 49 0 110 jjr ics=350uA

R0 VBIAS 41 80
R1 VBIAS 44 80
R2 VBIAS 49 40

RS0 40 41 3.9
RS1 41 0 3.9
RS2 43 0 2.7
RS3 42 43 3.9
RS4 47 49 3.9
RS5 50 44 3.9
RS6 44 0 3.9
RS7 46 0 2.7
RS8 45 46 3.9
RS9 48 49 3.9
RS10 49 0 1.9
.ends cin


.model jjr jj(level=2)
.tran 1p 0.8n
