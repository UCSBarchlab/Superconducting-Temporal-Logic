#! Delay Function Accelerator

* Testbench
.tran 1p 0.5n
.options ysep

.control
set Timestep=50p

set aVal=50p
*case 3 OK: 150p
*case 2 OK: 100p
*case 1 OK: 50p

set bVal=100p
*case 3: 150p
*case 2: 50p
*case 1: 100p

set cVal=150p
*case 3: 50p
*case 2: 5n
*case 1: 150p
.endc

V0 VCC 0 pwl 0 0 10p 10m


* Input Logic Pulses
Va 1 0 pulse 0 50m $aVal 50p 50p 100p 800p
Vb 3 0 pulse 0 50m $bVal 50p 50p 100p 800p
Vc 5 0 pulse 0 50m $cVal 50p 50p 100p 800p
* hard-coded '2' for second parameter set in table
Vh VTO 0 pulse 0 50m 100p 50p 50p 100p 800p
Vn VNM 0 pulse 0 0m 0p 50p 50p 100p 4n

* Input resistors
Ra 1 2 100
Rb 3 4 100
Rc 5 6 100
Rt VTO 8 100




* Macroscopic Delay Function

* Convert input pulses to SFQ
X0 2 IN1 VCC dcsfq
X1 4 IN2 VCC dcsfq
X2 6 IN3 VCC dcsfq
Xh 8 TWO VCC dcsfq

* Split each at first stage
X3 IN1 MD1s1 MD1s2 VCC split
X4 IN2 MD2s1 MD2s2 VCC split
X5 IN3 MD3s1 MD3s2 VCC split



* input to 1st logic block
* delay A = 150ps. Use "step" subckt, i.e. to make one time-step (50ps) worth of a delay
X6 MD1s1 MD1s11 VCC step
X7 MD1s11 MD1s12 VCC step
X8 MD1s12 MD1s13 VCC step
* B = 100ps
X15 MD2s1 MD2s11 VCC step
X16 MD2s11 MD2s12 VCC step
* C = 50ps
X20 MD3s1 MD3s11 VCC step

* 1st logic block 
X100 MD1s13 MD2s12 MD3s11 OUT1 VCC dfn





* input to 2nd logic block
X101 MD1s2 MD1s2s1 MD1s2s2 VCC split
X102 MD2s2 MD2s2s1 MD2s2s2 VCC split
X103 MD3s2 MD3s2s1 MD3s2s2 VCC split

X104 MD1s2s1 MD1211 VCC step
X105 MD2s2s1 MD2211 VCC step
X106 MD2211 MD2212 VCC step
X107 MD3s2s1 TWO MD3211 VCC inv
X108 MD3211 MD3212 VCC step2

* 2nd logic block
X200 MD1211 MD2212 MD3212 OUT2 VCC dfn



* input to 3rd logic block
X291 MD3s2s2 MD3221 VCC step
X292 MD3221 MD3222 VCC step

* 3rd logic block
X300 MD1s2s2 MD2s2s2 MD3222 OUT3 VCC dfn


*X414 COIN3 OUT3 VCC jtl


* First arrival
X301 OUT2 OUT3 OUT23 VCC merge
*X302 OUT1 OUT11 VCC jtl
*X303 OUT11 OUT12 VCC jtl
X304 OUT23 OUT1 FIRST VCC merge



* End of macroscopic Delay Function


* RSFQ Pulse Generation
.subckt dcsfq IN OUT VBIAS
B0 9 5 15 jjr ics=170uA
RS0 9 5 4
B1 10 11 16 jjr ics=250uA
RS1 10 11 2.7
B2 12 13 17 jjr ics=150uA
RS2 12 13 4.6
B3 7 14 18 jjr ics=170uA
RS3 7 14 4

L0 12 0 3.58pH
LP0 8 6 0.08pH
LP1 4 9 1.29pH
LP2 5 6 1.13pH
LP3 6 10 1.74pH
LP4 5 7 0.21pH
LP5 4 12 1.27pH
LP6 11 0 0.13pH
LP7 13 7 0.69pH
LP8 14 0 0.18pH

LT0 10 OUT 2.11pH
LT1 IN 4 3.38pH

R0 VBIAS 8 27
.ends dcsfq



* Delay function logic block for functions 1 and 2
.subckt dfn IN1 IN2 IN3 OUT VBIAS

X0 IN1 OUT11 OUT12 VBIAS split
X1 IN2 OUT21 OUT22 VBIAS split

* path balancing on 'c' line
X30 IN3 IN31 VBIAS jtl
X31 IN31 IN32 VBIAS jtl
X32 IN32 IN33 VBIAS jtl
X33 IN33 IN34 VBIAS jtl
X34 IN34 IN35 VBIAS jtl
X2 IN35 OUT31 OUT32 VBIAS split

X3 OUT11 OUT21 MERGE12 VBIAS merge
X4 MERGE12 MERGE121 VBIAS jtl
X5 MERGE121 MERGE122 VBIAS jtl

X6 OUT12 OUT22 MERGE122 COIN12 VBIAS cin

X7 COIN12 COIN1 COIN2 VBIAS split

X8 COIN1 OUT32 MERGE3 VBIAS merge
X409 MERGE3 MERGE31 VBIAS jtl
X410 MERGE31 MERGE32 VBIAS jtl
X13 COIN2 OUT31 MERGE32 COIN3 VBIAS cin

X14 COIN3 OUT VBIAS jtl

.ends dfn


* Splitter Element
.subckt split IN OUT1 OUT2 VBIAS
B0 2 0 100 jjr ics=355uA
R0 2 0 1.9
B1 7 0 101 jjr ics=250uA
R2 7 0 2.7
B2 9 0 102 jjr ics=250uA
R3 9 0 2.7

L0 IN 1 0.8p
L1 1 3 1.2p
L2 3 5 0.05p
L3 5 6 1.6p
L4 6 OUT1 1.98p
L5 5 8 1.6p
L6 8 OUT2 1.98p

LP0 1 2 0.05p
LP1 4 3 0.13p
LP2 6 7 0.05p
LP3 8 9 0.05p

R1 VBIAS 4 16.7
.ends split



* Merge Element
.subckt merge IN1 IN2 OUT VBIAS
B0 6 7 16 jjr ics=250uA
RS0 6 7 2.7
B1 8 10 17 jjr ics=224uA
RS1 8 10 3.4
B2 10 12 18 jjr ics=224uA
RS2 10 12 3.4
B3 11 13 19 jjr ics=250uA
RS3 11 13 2.7
B4 14 15 20 jjr ics=250uA
RS4 14 15 2.7

L0 IN1 7 6pH
L1 5 11 2.6pH
L2 11 OUT 2pH
L3 IN2 14 6pH

LP0 0 6 .03pH
LP1 7 8 .66pH
LP2 9 5 .13pH
LP3 10 5 .2pH
LP4 12 14 .66pH
LP5 13 0 .03pH
LP6 15 0 .03pH

R0 VBIAS 9 20
.ends merge


* Single Coincidence Element
.subckt cin IN1 IN2 CLK OUT VBIAS

* Clock signal is 
X5 CLK CLK1 CLK2 VBIAS split

L0 IN1 40 2p
L1 41 43 10p
L2 CLK1 42 2p
L3 43 47 4p
L4 IN2 50 2p
L5 44 46 10p
L6 CLK2 45 2p
L7 46 48 4p
L8 49 OUT 1.5p

B0 40 41 100 jjr ics=175uA
B1 41 0 101 jjr ics=175uA
B2 43 0 102 jjr ics=250uA
B3 42 43 103 jjr ics=175uA
B4 47 49 104 jjr ics=175uA
B5 50 44 105 jjr ics=175uA
B6 44 0 106 jjr ics=175uA
B7 46 0 107 jjr ics=250uA
B8 45 46 108 jjr ics=175uA
B9 48 49 109 jjr ics=175uA
B10 49 0 110 jjr ics=350uA

R0 VBIAS 41 80
R1 VBIAS 44 80
R2 VBIAS 49 40

RS0 40 41 3.9
RS1 41 0 3.9
RS2 43 0 2.7
RS3 42 43 3.9
RS4 47 49 3.9
RS5 50 44 3.9
RS6 44 0 3.9
RS7 46 0 2.7
RS8 45 46 3.9
RS9 48 49 3.9
RS10 49 0 1.9
.ends cin


* Inverter Element
.subckt inv 26 27 28 VBIAS
B0 10 11 29 jjr ics=140uA
RS0 10 11 4.9
B1 9 15 30 jjr ics=250uA
RS1 9 15 3.7
B2 10 16 31 jjr ics=310uA
RS2 10 16 2.2
B3 12 17 32 jjr ics=174uA
RS3 12 17 3.9
B4 13 18 33 jjr ics=294uA
RS4 13 18 2.3
B5 14 19 34 jjr ics=355uA
RS5 14 19 1.9
B6 21 24 35 jjr ics=294uA
RS6 21 24 2.3
B7 23 25 36 jjr ics=264uA
RS7 23 25 2.6

L0 26 9 2pH
L1 9 6 1.03pH
L2 6 10 .97pH
L3 11 12 .97pH
L4 12 7 .33pH
L5 7 13 5.88pH
L6 8 13 1.3pH
L7 14 8 1.02pH
L8 27 14 .79pH
L9 17 20 1.04pH
L10 20 18 .57pH
L11 20 21 .875pH
L12 21 22 1.7pH
L13 22 23 1.11pH
L14 23 28 2.37pH

LP0 3 6 .35pH
LP1 4 7 .57pH
LP2 5 8 .33pH
LP3 15 0 .03pH
LP4 16 0 .09pH
LP5 19 0 .02pH
LP6 2 22 .5pH
LP7 24 0 .145pH
LP8 25 0 .03pH

R0 VBIAS 3 40
R1 VBIAS 4 42
R2 VBIAS 5 74
R3 VBIAS 2 65
.ends inv



* Single JTL Circuit Element
.subckt jtl IN OUT VBIAS
B0 5 7 9 jjr ics=250uA
RS0 5 7 2.7
B1 6 8 10 jjr ics=250uA
RS1 6 8 2.7
LP0 7 0 .1pH
LP1 8 0 .1pH
LT0 IN 5 2.1pH
LT1 5 4 2.1pH
LT2 4 6 2.1pH
LT3 6 OUT 2.1pH
R0 VBIAS 4 29
.ends jtl


* Single delay time step (~50ps equivalent)
.subckt step IN OUT VBIAS
X0 IN 1 VBIAS jtl
X1 1 2 VBIAS jtl
X2 2 3 VBIAS jtl
X3 3 4 VBIAS jtl
X4 4 5 VBIAS jtl
X5 5 6 VBIAS jtl
X6 6 7 VBIAS jtl
X7 7 8 VBIAS jtl
X8 8 9 VBIAS jtl
X9 9 OUT VBIAS jtl
.ends step


* Single delay time step minus overhead of inverter in case 2 (~40ps equivalent)
.subckt step2 IN OUT VBIAS
X0 IN 1 VBIAS jtl
X1 1 2 VBIAS jtl
X2 2 3 VBIAS jtl
X3 3 4 VBIAS jtl
X4 4 5 VBIAS jtl
X5 5 6 VBIAS jtl
X6 6 7 VBIAS jtl
X7 7 8 VBIAS jtl
X8 8 OUT VBIAS jtl
.ends step2



.subckt buf IN OUT VBIAS
B0 2 0 100 jjr ics=355uA
RS0 2 0 1.9
B1 2 3 101 jjr ics=250uA
RS1 2 3 2.7

L1 IN 2 2p
L2 3 OUT 2p

R0 VBIAS 3 57
.ends buf


* Model Definition
.model jjr jj(level=2)
