#! First Arrival -- stateless

* In our temporal logic (under the assumption that shorter delays represent smaller values), First Arrival circuit realizes MIN function.

* For its stateless implementation, all needed is a Merge element.

* In contrast to its stateful version, the existing implementation generates multiple output events, which "violates" one of the main 
* Race Logic constraints for at most one event per "wire". In some cases though, such a relaxation may not cause any malfunction and lead
* to significant area and speed improvements.

.options ysep
R0 10 11 100
R1 20 21 100
V0 VCC 0 pwl 0 0 10p 10m

* Input Logic Pulses
V1 10 0 pulse 0 50m 50p 50p 50p 100p 350p
V2 20 0 pulse 0 50m 90p 50p 50p 20p 310p

* Macroscopic Stateless-First Arrival Circuit
X0 11 12 VCC dcsfq
X1 12 IN1 VCC jtl
X2 21 22 VCC dcsfq
X3 22 IN2 VCC jtl
X4 IN1 IN2 OUT VCC merge

* RSFQ Pulse Generation
* RS = JJ damping shunts, using Stewart-McCumber parameter with B_c = 1
.subckt dcsfq IN OUT VBIAS
B0 9 5 15 jjr ics=170uA
RS0 9 5 4
B1 10 11 16 jjr ics=250uA
RS1 10 11 2.7
B2 12 13 17 jjr ics=150uA
RS2 12 13 4.6
B3 7 14 18 jjr ics=170uA
RS3 7 14 4

L0 12 0 3.58pH
LP0 8 6 0.08pH
LP1 4 9 1.29pH
LP2 5 6 1.13pH
LP3 6 10 1.74pH
LP4 5 7 0.21pH
LP5 4 12 1.27pH
LP6 11 0 0.13pH
LP7 13 7 0.69pH
LP8 14 0 0.18pH

LT0 10 OUT 2.11pH
LT1 IN 4 3.38pH

R0 VBIAS 8 27
.ends dcsfq

* Single JTL Circuit Element
.subckt jtl IN OUT VBIAS
B0 5 7 9 jjr ics=250uA
RS0 5 7 2.7
B1 6 8 10 jjr ics=250uA
RS1 6 8 2.7

LP0 7 0 .1pH
LP1 8 0 .1pH

LT0 IN 5 2.1pH
LT1 5 4 2.1pH
LT2 4 6 2.1pH
LT3 6 OUT 2.1pH

R0 VBIAS 4 29
.ends jtl

* Merge Element
.subckt merge IN1 IN2 OUT VBIAS
B0 6 7 16 jjr ics=250uA
RS0 6 7 2.7
B1 8 10 17 jjr ics=220uA
RS1 8 10 3.1
B2 10 12 18 jjr ics=220uA
RS2 10 12 3.1
B3 11 13 19 jjr ics=250uA
RS3 11 13 2.7
B4 14 15 20 jjr ics=250uA
RS4 14 15 2.7

L0 IN1 7 5pH
L1 5 11 2.6pH
L2 11 OUT 2pH
L3 IN2 14 5pH

LP0 0 6 .03pH
LP1 7 8 .66pH
LP2 9 5 .13pH
LP3 10 5 .2pH
LP4 12 14 .66pH
LP5 13 0 .03pH
LP6 15 0 .03pH

R0 VBIAS 9 20
.ends merge

* Model Definition
.model jjr jj(level=2)

.tran 1p 0.6n
